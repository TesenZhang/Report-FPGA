module vga_pic(
input wire vga_clk , 
input wire sys_rst_n , 
input wire [9:0] pix_x , 
input wire [9:0] pix_y , 

output reg [15:0] pix_data 

);


parameter CHAR_B_H= 10'd192 , 
CHAR_B_V= 10'd208 ; 

parameter CHAR_W = 10'd256 , 
CHAR_H = 10'd64 ; 

parameter BLACK = 16'h0000, 
WHITE = 16'hFFFF, 
GOLDEN = 16'hFEC0; 


wire [9:0] char_x ; 
wire [9:0] char_y ; 


reg [255:0] char [63:0] ; 
assign char_x=(((pix_x>=CHAR_B_H) && (pix_y<(CHAR_B_H+CHAR_W)))
					&&((pix_y>=CHAR_B_V) &&(pix_y<(CHAR_B_V+CHAR_H)) ))
					? (pix_x - CHAR_B_H) :10'h3ff;
assign char_y = (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
&&((pix_y >= CHAR_B_V)&&(pix_y < (CHAR_B_V + CHAR_H))))
? (pix_y - CHAR_B_V) : 10'h3FF;
					


always@(posedge vga_clk)
    begin
        char[0]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[1]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[2]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[3]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[4]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[5]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[6]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[7]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[8]  <= 256'h0000000000000000000000000000000000000000000000000003FC0000000000;
        char[9]  <= 256'h3F8000FE3E00007E003FFFF07FFFFFFF3F8001FE3E00007E00FFFFF07FFFFFFF;
        char[10] <= 256'h3FC001FE3E00007E03FFFFF07FFFFFFF3FC001FE3E00007E07FFFFF07FFFFFFF;
        char[11] <= 256'h7FC003FE3E00007E0FF800F00007E0007FE003FE3E00007E1FE000000007E000;
        char[12] <= 256'h7FE007FF3E00007E1F8000000007E0007DF007FF3E00007E1F8000000007E000;
        char[13] <= 256'h7DF007BF3E00007E3F0000000007E0007DF00FBF3E00007E3F0000000007E000;
        char[14] <= 256'h7CF80F1F3E00007E3F0000000007E0007CF81F1F3E00007E3F8000000007E000;
        char[15] <= 256'h7CF81F1F3E00007E3F8000000007E0007C7C1E1F3E00007E1FC000000007E000;
        char[16] <= 256'h7C7C3E1F3E00007E1FE000000007E0007C3E3E1F3E00007E0FF800000007E000;
        char[17] <= 256'h7C3E7C1F3E00007E07FF00000007E0007C3E7C1F3E00007E03FFC0000007E000;
        char[18] <= 256'h7C1F781F3E00007E01FFF8000007E0007C1FF81F3E00007E007FFE000007E000;
        char[19] <= 256'h7C1FF81F3E00007E001FFF800007E0007C0FF01F3E00007E0003FFE00007E000;
        char[20] <= 256'h7C0FF01F3E00007E0000FFF00007E000FC07E01F3E00007E00001FF80007E000;
        char[21] <= 256'hFC07E01F3E00007E000007F80007E000FC07E01F3E00007E000003FC0007E000;
        char[22] <= 256'hFC03C01F3E00007E000001FC0007E000F800001F3E00007E000000FC0007E000;
        char[23] <= 256'hF800001F3E00007E000000FE0007E000F800001F3F00007E0000007E0007E000;
        char[24] <= 256'hF800001F3F00007E000000FE0007E000F800001F3F00007C000000FC0007E000;
        char[25] <= 256'hF800001F3F8000FC000000FC0007E000F800001F1F8001FC000001FC0007E000;
        char[26] <= 256'hF800001F1FE003F8300007F80007E000F800001F0FF80FF03F803FF00007E000;
        char[27] <= 256'hF800001F07FFFFE03FFFFFE00007E000F800001F03FFFFC03FFFFFC00007E000;
        char[28] <= 256'hF800001F01FFFF803FFFFF000007E000F800000F007FFE001FFFFC000007E000;
        char[29] <= 256'h000000000001C000000F00000000000000000000000000000000000000000000;
        char[30] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[31] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[32] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[33] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[34] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[35] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[36] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[37] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[38] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[39] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[40] <= 256'h0000000000000000000000000000000000000000000000000003FC0000000000;
        char[41] <= 256'h3F8000FE3E00007E003FFFF07FFFFFFF3F8001FE3E00007E00FFFFF07FFFFFFF;
        char[42] <= 256'h3FC001FE3E00007E03FFFFF07FFFFFFF3FC001FE3E00007E07FFFFF07FFFFFFF;
        char[43] <= 256'h7FC003FE3E00007E0FF800F00007E0007FE003FE3E00007E1FE000000007E000;
        char[44] <= 256'h7FE007FF3E00007E1F8000000007E0007DF007FF3E00007E1F8000000007E000;
        char[45] <= 256'h7DF007BF3E00007E3F0000000007E0007DF00FBF3E00007E3F0000000007E000;
        char[46] <= 256'h7CF80F1F3E00007E3F0000000007E0007CF81F1F3E00007E3F8000000007E000;
        char[47] <= 256'h7CF81F1F3E00007E3F8000000007E0007C7C1E1F3E00007E1FC000000007E000;
        char[48] <= 256'h7C7C3E1F3E00007E1FE000000007E0007C3E3E1F3E00007E0FF800000007E000;
        char[49] <= 256'h7C3E7C1F3E00007E07FF00000007E0007C3E7C1F3E00007E03FFC0000007E000;
        char[50] <= 256'h7C1F781F3E00007E01FFF8000007E0007C1FF81F3E00007E007FFE000007E000;
        char[51] <= 256'h7C1FF81F3E00007E001FFF800007E0007C0FF01F3E00007E0003FFE00007E000;
        char[52] <= 256'h7C0FF01F3E00007E0000FFF00007E000FC07E01F3E00007E00001FF80007E000;
        char[53] <= 256'hFC07E01F3E00007E000007F80007E000FC07E01F3E00007E000003FC0007E000;
        char[54] <= 256'hFC03C01F3E00007E000001FC0007E000F800001F3E00007E000000FC0007E000;
        char[55] <= 256'hF800001F3E00007E000000FE0007E000F800001F3F00007E0000007E0007E000;
        char[56] <= 256'hF800001F3F00007E000000FE0007E000F800001F3F00007C000000FC0007E000;
        char[57] <= 256'hF800001F3F8000FC000000FC0007E000F800001F1F8001FC000001FC0007E000;
        char[58] <= 256'hF800001F1FE003F8300007F80007E000F800001F0FF80FF03F803FF00007E000;
        char[59] <= 256'hF800001F07FFFFE03FFFFFE00007E000F800001F03FFFFC03FFFFFC00007E000;
        char[60] <= 256'hF800001F01FFFF803FFFFF000007E000F800000F007FFE001FFFFC000007E000;
        char[61] <= 256'h000000000001C000000F00000000000000000000000000000000000000000000;
        char[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    end                  
	 
 always@(posedge vga_clk or negedge sys_rst_n)
 if(sys_rst_n == 1'b0)
 pix_data <= BLACK;
 else if((((pix_x >= (CHAR_B_H - 1'b1))
 && (pix_x < (CHAR_B_H + CHAR_W -1'b1)))
 && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
 && (char[char_y][10'd255 - char_x] == 1'b1))
 pix_data <= GOLDEN;
 else
 pix_data <= BLACK;

 endmodule